    x"7e517e51",
    x"87408740",
    x"90409040",
    x"137f137f",
    x"3d0d3d0d",
    x"500a500a",
    x"d668d668",
    x"b1d7b1d7",
    x"44694469",
    x"dd06dd06",
    x"bcaabcaa",
    x"1ea81ea8",
    x"97ae97ae",
    x"cd45cd45",
    x"2d2d2d2d",
    x"b5a1b5a1",
    x"b307b307",
    x"9fb39fb3",
    x"91179117",
    x"93429342",
    x"18261826",
    x"78bd78bd",
    x"ba00ba00",
    x"53e053e0",
    x"077c077c",
    x"201f201f",
    x"bb40bb40",
    x"cbb9cbb9",
    x"37083708",
    x"29852985",
    x"eef3eef3",
    x"b55ab55a",
    x"b0c5b0c5",
    x"7f337f33",
    x"c8d9c8d9",
    x"edd2edd2",
    x"cf3dcf3d",
    x"9f419f41",
    x"9fa99fa9",
    x"13a713a7",
    x"7c487c48",
    x"5c535c53",
    x"324f324f",
    x"13f613f6",
    x"29992999",
    x"5f7d5f7d",
    x"c997c997",
    x"dca0dca0",
    x"ff30ff30",
    x"5aae5aae",
    x"6fe36fe3",
    x"17561756",
    x"d36bd36b",
    x"29e329e3",
    x"6b376b37",
    x"dae7dae7",
    x"4a024a02",
    x"26772677",
    x"a6a1a6a1",
    x"810b810b",
    x"4ffc4ffc",
    x"95949594",
    x"36653665",
    x"00c100c1"